module ALU(

	input 	wire[15:0] 	wInstruction;
	

);
